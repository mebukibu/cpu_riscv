`include "consts.vh"

// load, store
`define LW      `WORD_LEN'b00000000000000000010000000000011     // type I
`define SW      `WORD_LEN'b00000000000000000010000000100011     // type S

// add
`define ADD     `WORD_LEN'b00000000000000000000000000110011     // type R
`define ADDI    `WORD_LEN'b00000000000000000000000000010011     // type I

// sub
`define SUB     `WORD_LEN'b01000000000000000000000000110011     // type R

// logic
`define AND     `WORD_LEN'b00000000000000000111000000110011     // type R
`define OR      `WORD_LEN'b00000000000000000110000000110011     // type R
`define XOR     `WORD_LEN'b00000000000000000100000000110011     // type R
`define ANDI    `WORD_LEN'b00000000000000000111000000010011     // type I
`define ORI     `WORD_LEN'b00000000000000000110000000010011     // type I
`define XORI    `WORD_LEN'b00000000000000000100000000010011     // type I

// shift
`define SLL     `WORD_LEN'b0000000XXXXXXXXXX001XXXXX0110011
`define SRL     `WORD_LEN'b0000000XXXXXXXXXX101XXXXX0110011
`define SRA     `WORD_LEN'b0100000XXXXXXXXXX101XXXXX0110011
`define SLLI    `WORD_LEN'b0000000XXXXXXXXXX001XXXXX0010011
`define SRLI    `WORD_LEN'b0000000XXXXXXXXXX101XXXXX0010011
`define SRAI    `WORD_LEN'b0100000XXXXXXXXXX101XXXXX0010011

// comparison
`define SLT     `WORD_LEN'b0000000XXXXXXXXXX010XXXXX0110011
`define SLTU    `WORD_LEN'b0000000XXXXXXXXXX011XXXXX0110011
`define SLTI    `WORD_LEN'bXXXXXXXXXXXXXXXXX010XXXXX0010011
`define SLTIU   `WORD_LEN'bXXXXXXXXXXXXXXXXX011XXXXX0010011

// conditional branch
`define BEQ     `WORD_LEN'bXXXXXXXXXXXXXXXXX000XXXXX1100011
`define BNE     `WORD_LEN'bXXXXXXXXXXXXXXXXX001XXXXX1100011
`define BLT     `WORD_LEN'bXXXXXXXXXXXXXXXXX100XXXXX1100011
`define BGE     `WORD_LEN'bXXXXXXXXXXXXXXXXX101XXXXX1100011
`define BLTU    `WORD_LEN'bXXXXXXXXXXXXXXXXX110XXXXX1100011
`define BGEU    `WORD_LEN'bXXXXXXXXXXXXXXXXX111XXXXX1100011

// jump
`define JAL     `WORD_LEN'bXXXXXXXXXXXXXXXXXXXXXXXXX1101111
`define JALR    `WORD_LEN'bXXXXXXXXXXXXXXXXX000XXXXX1100111

// im load
`define LUI     `WORD_LEN'bXXXXXXXXXXXXXXXXXXXXXXXXX0110111
`define AUIPC   `WORD_LEN'bXXXXXXXXXXXXXXXXXXXXXXXXX0010111

// CSR
`define CSRRW   `WORD_LEN'bXXXXXXXXXXXXXXXXX001XXXXX1110011
`define CSRRWI  `WORD_LEN'bXXXXXXXXXXXXXXXXX101XXXXX1110011
`define CSRRS   `WORD_LEN'bXXXXXXXXXXXXXXXXX010XXXXX1110011
`define CSRRSI  `WORD_LEN'bXXXXXXXXXXXXXXXXX110XXXXX1110011
`define CSRRC   `WORD_LEN'bXXXXXXXXXXXXXXXXX011XXXXX1110011
`define CSRRCI  `WORD_LEN'bXXXXXXXXXXXXXXXXX111XXXXX1110011

// except
`define ECALL   `WORD_LEN'b00000000000000000000000001110011

// vector
`define VSETVLI `WORD_LEN'bXXXXXXXXXXXXXXXXX111XXXXX1010111
`define VLE     `WORD_LEN'b000000100000XXXXXXXXXXXXX0000111
`define VSE     `WORD_LEN'b000000100000XXXXXXXXXXXXX0100111
`define VADDVV  `WORD_LEN'b0000001XXXXXXXXXX000XXXXX1010111

// custom
`define PCNT    `WORD_LEN'b000000000000XXXXX110XXXXX0001011


// instruction type mask
`define TYPE_R  `WORD_LEN'b11111110000000000111000001111111
`define TYPE_IS `WORD_LEN'b00000000000000000111000001111111
`define TYPE_U  `WORD_LEN'b00000000000000000000000001111111